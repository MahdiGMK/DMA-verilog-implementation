module dma ();

endmodule
