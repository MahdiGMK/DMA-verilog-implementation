module cpu ();
endmodule
